//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company : AGH University of Krakow
// Create Date : 23.07.2024
// Designers Name : Dawid Mironiuk & Michał Malara
// Module Name : figure_rom
// Project Name : SZACHY - Projekt zaliczeniowy
// Target Devices : BASYS3
// 
// Description : Moduł odpowiedzialny za wygląd czcionki figur.
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module figure_rom
    (
        input  logic        clk,
        input  logic [8:0] addr,                 // {figure_code[5:0], figure_line[4:0]} //
        output logic  [63:0] figure_line_pixels   // pixels of the figure line //
    );

    // SIGNAL DECLARATION //////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

    logic [63:0] data;

    // BODY ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

    always_ff @(posedge clk) begin
        //figure_line_pixels <= data;
    //end
        
    //always_comb begin
        case (addr)
            // 00-bg 01-szary 10-biła 11-czarny
            // CODE x00 PUSTE POLE //////////////
            9'h000: data <= 64'h0000000000000000;
            9'h001: data <= 64'h0000000000000000;
            9'h002: data <= 64'h0000000000000000;
            9'h003: data <= 64'h0000000000000000;
            9'h004: data <= 64'h0000000000000000;
            9'h005: data <= 64'h0000000000000000;
            9'h006: data <= 64'h0000000000000000;
            9'h007: data <= 64'h0000000000000000;
            9'h008: data <= 64'h0000000000000000;
            9'h009: data <= 64'h0000000000000000;
            9'h00a: data <= 64'h0000000000000000;
            9'h00b: data <= 64'h0000000000000000;
            9'h00c: data <= 64'h0000000000000000;
            9'h00d: data <= 64'h0000000000000000;
            9'h00e: data <= 64'h0000000000000000;
            9'h00f: data <= 64'h0000000000000000;
            9'h010: data <= 64'h0000000000000000;
            9'h011: data <= 64'h0000000000000000;
            9'h012: data <= 64'h0000000000000000;
            9'h013: data <= 64'h0000000000000000;
            9'h014: data <= 64'h0000000000000000;
            9'h015: data <= 64'h0000000000000000;
            9'h016: data <= 64'h0000000000000000;
            9'h017: data <= 64'h0000000000000000;
            9'h018: data <= 64'h0000000000000000;
            9'h019: data <= 64'h0000000000000000;
            9'h01a: data <= 64'h0000000000000000;
            9'h01b: data <= 64'h0000000000000000; 
            9'h01c: data <= 64'h0000000000000000;
            9'h01d: data <= 64'h0000000000000000;
            9'h01e: data <= 64'h0000000000000000;
            9'h01f: data <= 64'h0000000000000000;
            // CODE x01 BIAŁY PIONEK ////////////
            9'h020: data <= 64'h0000000000000000; 
            9'h021: data <= 64'h0000000000000000;
            9'h022: data <= 64'h0000000000000000;
            9'h023: data <= 64'h0000000000000000;
            9'h024: data <= 64'h0000000000000000;
            9'h025: data <= 64'h0000000000000000;
            9'h026: data <= 64'h0000000000000000;
            9'h027: data <= 64'h0000000000000000;
            9'h028: data <= 64'h0000000000000000;
            9'h029: data <= 64'h0000000000000000;
            9'h02a: data <= 64'h0000000000000000;
            9'h02b: data <= 64'h0000000000000000;
            9'h02c: data <= 64'h0000000550000000;
            9'h02d: data <= 64'h0000001AA4000000;
            9'h02e: data <= 64'h0000006AA9000000;
            9'h02f: data <= 64'h0000006AA9000000;
            9'h030: data <= 64'h0000006AA9000000;
            9'h031: data <= 64'h0000006AA9000000;
            9'h032: data <= 64'h0000001AA4000000;
            9'h033: data <= 64'h0000000690000000;
            9'h034: data <= 64'h0000000690000000;
            9'h035: data <= 64'h0000001AA4000000;
            9'h036: data <= 64'h0000001AA4000000;
            9'h037: data <= 64'h0000006AA9000000;
            9'h038: data <= 64'h0000006AA9000000;
            9'h039: data <= 64'h000001AAAA400000;
            9'h03a: data <= 64'h000001AAAA400000;
            9'h03b: data <= 64'h0000055555500000;
            9'h03c: data <= 64'h000006AAAA900000;
            9'h03d: data <= 64'h0000055555500000;
            9'h03e: data <= 64'h0000000000000000;
            9'h03f: data <= 64'h0000000000000000;
            // CODE x02 BIAŁY GONIEC //////////// 
            9'h040: data <= 64'h0000000000000000;
            9'h041: data <= 64'h0000000000000000;
            9'h042: data <= 64'h0000000140000000;
            9'h043: data <= 64'h0000000690000000;
            9'h044: data <= 64'h0000000690000000;
            9'h045: data <= 64'h0000000140000000;
            9'h046: data <= 64'h0000000690000000;
            9'h047: data <= 64'h0000001AA4000000;
            9'h048: data <= 64'h0000006AA9000000;
            9'h049: data <= 64'h000001AAAA400000;
            9'h04a: data <= 64'h000001AAAA400000;
            9'h04b: data <= 64'h000006AAA9000000;
            9'h04c: data <= 64'h00001AAAA4140000;
            9'h04d: data <= 64'h00001AAA90640000;
            9'h04e: data <= 64'h00006AAA91A90000;
            9'h04f: data <= 64'h00006AAAA6A90000;
            9'h050: data <= 64'h00006AAAAAA90000;
            9'h051: data <= 64'h00006AAAAAA90000;
            9'h052: data <= 64'h00001AAAAAA40000;
            9'h053: data <= 64'h00001AAAAAA40000;
            9'h054: data <= 64'h00001AAAAAA40000;
            9'h055: data <= 64'h000006AAAA900000;
            9'h056: data <= 64'h000006AAAA900000;
            9'h057: data <= 64'h000001AAAA400000;
            9'h058: data <= 64'h000001AAAA400000;
            9'h059: data <= 64'h0000055555500000;
            9'h05a: data <= 64'h00001AAAAAA40000;
            9'h05b: data <= 64'h0000555555550000;
            9'h05c: data <= 64'h00006AAAAAA90000;
            9'h05d: data <= 64'h0000555555550000;
            9'h05e: data <= 64'h0000000000000000;
            9'h05f: data <= 64'h0000000000000000;
            // CODE x03 BIAŁY KOŃ ///////////////
            9'h060: data <= 64'h0000000000000000;
            9'h061: data <= 64'h0000000000000000;
            9'h062: data <= 64'h0000000000000000;
            9'h063: data <= 64'h0000000000000000;
            9'h064: data <= 64'h0000000000000000;
            9'h065: data <= 64'h0000000000000000;
            9'h066: data <= 64'h0000000000000000;
            9'h067: data <= 64'h0000005400000000;
            9'h068: data <= 64'h000001A954000000;
            9'h069: data <= 64'h000001AAA9400000;
            9'h06a: data <= 64'h0000005AAA900000;
            9'h06b: data <= 64'h00000006AAA40000;
            9'h06c: data <= 64'h0000001AAAA50000;
            9'h06d: data <= 64'h00000169AAA90000;
            9'h06e: data <= 64'h000006AAAAA90000;
            9'h06f: data <= 64'h000006AAAAA90000;
            9'h070: data <= 64'h00001AAAAAA90000;
            9'h071: data <= 64'h00006AA5AAA90000;
            9'h072: data <= 64'h00006951AAA40000;
            9'h073: data <= 64'h00001401AAA40000;
            9'h074: data <= 64'h00000006AAA40000;
            9'h075: data <= 64'h0000001AAAA40000;
            9'h076: data <= 64'h0000006AAA900000;
            9'h077: data <= 64'h000001AAAA900000;
            9'h078: data <= 64'h000001AAAA900000;
            9'h079: data <= 64'h0000055555500000;
            9'h07a: data <= 64'h00001AAAAAA40000;
            9'h07b: data <= 64'h0000555555550000;
            9'h07c: data <= 64'h00006AAAAAA90000;
            9'h07d: data <= 64'h0000555555550000;
            9'h07e: data <= 64'h0000000000000000;
            9'h07f: data <= 64'h0000000000000000;
            // CODE x04 WIEŻA BIAŁA /////////////
            9'h080: data <= 64'h0000000000000000; 
            9'h081: data <= 64'h0000000000000000;
            9'h082: data <= 64'h0000000000000000;
            9'h083: data <= 64'h0000000000000000;
            9'h084: data <= 64'h0000000000000000;
            9'h085: data <= 64'h0000000000000000;
            9'h086: data <= 64'h0000000000000000;
            9'h087: data <= 64'h0000000000000000;
            9'h088: data <= 64'h0000551554550000;
            9'h089: data <= 64'h00006A5AA5A90000;
            9'h08a: data <= 64'h00006AAAAAA90000;
            9'h08b: data <= 64'h00005AAAAAA50000;
            9'h08c: data <= 64'h0000155555540000;
            9'h08d: data <= 64'h000006AAAA900000;
            9'h08e: data <= 64'h0000055555500000;
            9'h08f: data <= 64'h000001AAAA400000;
            9'h090: data <= 64'h000001AAAA400000;
            9'h091: data <= 64'h000001AAAA400000;
            9'h092: data <= 64'h000001AAAA400000;
            9'h093: data <= 64'h000001AAAA400000;
            9'h094: data <= 64'h000001AAAA400000;
            9'h095: data <= 64'h000001AAAA400000;
            9'h096: data <= 64'h000001AAAA400000;
            9'h097: data <= 64'h000001AAAA400000;
            9'h098: data <= 64'h0000055555500000;
            9'h099: data <= 64'h000006AAAA900000;
            9'h09a: data <= 64'h0000155555540000;
            9'h09b: data <= 64'h00005AAAAAA50000;
            9'h09c: data <= 64'h00006AAAAAA90000;
            9'h09d: data <= 64'h0000555555550000;
            9'h09e: data <= 64'h0000000000000000;
            9'h09f: data <= 64'h0000000000000000;
            // CODE x05 KRÓLOWA BIAŁA ///////////
            9'h0a0: data <= 64'h0000000000000000; 
            9'h0a1: data <= 64'h0000000000000000;
            9'h0a2: data <= 64'h0000000000000000;
            9'h0a3: data <= 64'h0000000000000000;
            9'h0a4: data <= 64'h0000000000000000;
            9'h0a5: data <= 64'h0000000000000000;
            9'h0a6: data <= 64'h0000000000000000;
            9'h0a7: data <= 64'h0000000000000000;
            9'h0a8: data <= 64'h0000000000000000;
            9'h0a9: data <= 64'h0000000000000000;
            9'h0aa: data <= 64'h0000000000000000;
            9'h0ab: data <= 64'h0000000000000000;
            9'h0ac: data <= 64'h0001400140014000;
            9'h0ad: data <= 64'h0001900690064000;
            9'h0ae: data <= 64'h0001A406901A4000;
            9'h0af: data <= 64'h0001A901406A4000;
            9'h0b0: data <= 64'h0001A906906A4000;
            9'h0b1: data <= 64'h0001AA5AA5AA4000;
            9'h0b2: data <= 64'h0001AAAAAAAA4000;
            9'h0b3: data <= 64'h0001AAAAAAAA4000;
            9'h0b4: data <= 64'h00006AAAAAA90000;
            9'h0b5: data <= 64'h00001AAAAAA40000;
            9'h0b6: data <= 64'h0000055555500000;
            9'h0b7: data <= 64'h000006AAAA900000;
            9'h0b8: data <= 64'h000001AAAA400000;
            9'h0b9: data <= 64'h0000155555540000;
            9'h0ba: data <= 64'h00001AAAAAA40000;
            9'h0bb: data <= 64'h0000555555550000;
            9'h0bc: data <= 64'h00006AAAAAA90000;
            9'h0bd: data <= 64'h0000555555550000;
            9'h0be: data <= 64'h0000000000000000;
            9'h0bf: data <= 64'h0000000000000000;
            // CODE x06 KRÓL BIAŁY///////////////
            9'h0c0: data <= 64'h0000000000000000; 
            9'h0c1: data <= 64'h0000000000000000;
            9'h0c2: data <= 64'h0000000000000000;
            9'h0c3: data <= 64'h0000000000000000;
            9'h0c4: data <= 64'h0000000000000000;
            9'h0c5: data <= 64'h0000000000000000;
            9'h0c6: data <= 64'h0000000000000000;
            9'h0c7: data <= 64'h0000000140000000;
            9'h0c8: data <= 64'h0000000690000000;
            9'h0c9: data <= 64'h0000001694000000;
            9'h0ca: data <= 64'h0000006AA9000000;
            9'h0cb: data <= 64'h0000006AA9000000;
            9'h0cc: data <= 64'h0000001694000000;
            9'h0cd: data <= 64'h0000550690550000;
            9'h0ce: data <= 64'h0001AA5695AA4000;
            9'h0cf: data <= 64'h0006AAA69AAA9000;
            9'h0d0: data <= 64'h0006AAA96AAA9000;
            9'h0d1: data <= 64'h0006AAA96AAA9000;
            9'h0d2: data <= 64'h0006AAAAAAAA9000;
            9'h0d3: data <= 64'h0006AAAAAAAA9000;
            9'h0d4: data <= 64'h0006AAAAAAAA9000;
            9'h0d5: data <= 64'h0006AAAAAAAA9000;
            9'h0d6: data <= 64'h0001AAAAAAAA4000;
            9'h0d7: data <= 64'h0001AAAAAAAA4000;
            9'h0d8: data <= 64'h00006AAAAAA90000;
            9'h0d9: data <= 64'h0000155555540000;
            9'h0da: data <= 64'h00001AAAAAA40000;
            9'h0db: data <= 64'h0000555555550000;
            9'h0dc: data <= 64'h00006AAAAAA90000;
            9'h0dd: data <= 64'h0000555555550000;
            9'h0de: data <= 64'h0000000000000000;
            9'h0df: data <= 64'h0000000000000000;   
            // CODE x07 PIONEK CZARNY ///////////
            9'h0e0: data <= 64'h0000000000000000;   
            9'h0e1: data <= 64'h0000000000000000;
            9'h0e2: data <= 64'h0000000000000000;
            9'h0e3: data <= 64'h0000000000000000;
            9'h0e4: data <= 64'h0000000000000000;
            9'h0e5: data <= 64'h0000000000000000;
            9'h0e6: data <= 64'h0000000000000000;
            9'h0e7: data <= 64'h0000000000000000;
            9'h0e8: data <= 64'h0000000000000000;
            9'h0e9: data <= 64'h0000000000000000;
            9'h0ea: data <= 64'h0000000000000000;
            9'h0eb: data <= 64'h0000000000000000;
            9'h0ec: data <= 64'h0000000550000000;
            9'h0ed: data <= 64'h0000001FF4000000;
            9'h0ee: data <= 64'h0000007FFD000000;
            9'h0ef: data <= 64'h0000007FFD000000;
            9'h0f0: data <= 64'h0000007FFD000000;
            9'h0f1: data <= 64'h0000007FFD000000;
            9'h0f2: data <= 64'h0000001FF4000000;
            9'h0f3: data <= 64'h00000007D0000000;
            9'h0f4: data <= 64'h00000007D0000000;
            9'h0f5: data <= 64'h0000001FF4000000;
            9'h0f6: data <= 64'h0000001FF4000000;
            9'h0f7: data <= 64'h0000007FFD000000;
            9'h0f8: data <= 64'h0000007FFD000000;
            9'h0f9: data <= 64'h000001FFFF400000;
            9'h0fa: data <= 64'h000001FFFF400000;
            9'h0fb: data <= 64'h0000055555500000;
            9'h0fc: data <= 64'h000007FFFFD00000;
            9'h0fd: data <= 64'h0000055555500000;
            9'h0fe: data <= 64'h0000000000000000;
            9'h0ff: data <= 64'h0000000000000000;
            // CODE x08 GONIEC CZARNY ///////////
            9'h100: data <= 64'h0000000000000000;
            9'h101: data <= 64'h0000000000000000;
            9'h102: data <= 64'h0000000140000000;
            9'h103: data <= 64'h00000007D0000000;
            9'h104: data <= 64'h00000007D0000000;
            9'h105: data <= 64'h0000000140000000;
            9'h106: data <= 64'h00000007D0000000;
            9'h107: data <= 64'h0000001FF4000000;
            9'h108: data <= 64'h0000007FFD000000;
            9'h109: data <= 64'h000001FFFF400000;
            9'h10a: data <= 64'h000001FFFF400000;
            9'h10b: data <= 64'h000007FFFD000000;
            9'h10c: data <= 64'h00001FFFF4140000;
            9'h10d: data <= 64'h00001FFFD0740000;
            9'h10e: data <= 64'h00007FFFD1FD0000;
            9'h10f: data <= 64'h00007FFFF7FD0000;
            9'h110: data <= 64'h00007FFFFFFD0000;
            9'h111: data <= 64'h00007FFFFFFD0000;
            9'h112: data <= 64'h00001FFFFFF40000;
            9'h113: data <= 64'h00001FFFFFF40000;
            9'h114: data <= 64'h00001FFFFFF40000;
            9'h115: data <= 64'h000007FFFFD00000;
            9'h116: data <= 64'h000007FFFFD00000;
            9'h117: data <= 64'h000001FFFF400000;
            9'h118: data <= 64'h000001FFFF400000;
            9'h119: data <= 64'h0000055555500000;
            9'h11a: data <= 64'h00001FFFFFF40000;
            9'h11b: data <= 64'h0000555555550000;
            9'h11c: data <= 64'h00007FFFFFFD0000;
            9'h11d: data <= 64'h0000555555550000;
            9'h11e: data <= 64'h0000000000000000;
            9'h11f: data <= 64'h0000000000000000;
            // CODE x09 KOŃ CZARNY //////////////
            9'h120: data <= 64'h0000000000000000; 
            9'h121: data <= 64'h0000000000000000;
            9'h122: data <= 64'h0000000000000000;
            9'h123: data <= 64'h0000000000000000;
            9'h124: data <= 64'h0000000000000000;
            9'h125: data <= 64'h0000000000000000;
            9'h126: data <= 64'h0000000000000000;
            9'h127: data <= 64'h0000005400000000;
            9'h128: data <= 64'h000001FD54000000;
            9'h129: data <= 64'h000001FFFD400000;
            9'h12a: data <= 64'h0000005FFFD00000;
            9'h12b: data <= 64'h00000007FFF40000;
            9'h12c: data <= 64'h0000001FFFF50000;
            9'h12d: data <= 64'h0000017DFFFD0000;
            9'h12e: data <= 64'h000007FFFFFD0000;
            9'h12f: data <= 64'h000007FFFFFD0000;
            9'h130: data <= 64'h00001FFFFFFD0000;
            9'h131: data <= 64'h00007FF5FFFD0000;
            9'h132: data <= 64'h00007D51FFF40000;
            9'h133: data <= 64'h00001401FFF40000;
            9'h134: data <= 64'h00000007FFF40000;
            9'h135: data <= 64'h0000001FFFF40000;
            9'h136: data <= 64'h0000007FFFD00000;
            9'h137: data <= 64'h000001FFFFD00000;
            9'h138: data <= 64'h000001FFFFD00000;
            9'h139: data <= 64'h0000055555500000;
            9'h13a: data <= 64'h00001FFFFFF40000;
            9'h13b: data <= 64'h0000555555550000;
            9'h13c: data <= 64'h00007FFFFFFD0000;
            9'h13d: data <= 64'h0000555555550000;
            9'h13e: data <= 64'h0000000000000000;
            9'h13f: data <= 64'h0000000000000000;
            // CODE x10 WIEŻA CZARNA ////////////
            9'h140: data <= 64'h0000000000000000; 
            9'h141: data <= 64'h0000000000000000;
            9'h142: data <= 64'h0000000000000000;
            9'h143: data <= 64'h0000000000000000;
            9'h144: data <= 64'h0000000000000000;
            9'h145: data <= 64'h0000000000000000;
            9'h146: data <= 64'h0000000000000000;
            9'h147: data <= 64'h0000000000000000;
            9'h148: data <= 64'h0000551554550000;
            9'h149: data <= 64'h00007F5FF5FD0000;
            9'h14a: data <= 64'h00007FFFFFFD0000;
            9'h14b: data <= 64'h00005FFFFFF50000;
            9'h14c: data <= 64'h0000155555540000;
            9'h14d: data <= 64'h000007FFFFD00000;
            9'h14e: data <= 64'h0000055555500000;
            9'h14f: data <= 64'h000001FFFF400000;
            9'h150: data <= 64'h000001FFFF400000;
            9'h151: data <= 64'h000001FFFF400000;
            9'h152: data <= 64'h000001FFFF400000;
            9'h153: data <= 64'h000001FFFF400000;
            9'h154: data <= 64'h000001FFFF400000;
            9'h155: data <= 64'h000001FFFF400000;
            9'h156: data <= 64'h000001FFFF400000;
            9'h157: data <= 64'h000001FFFF400000;
            9'h158: data <= 64'h0000055555500000;
            9'h159: data <= 64'h000007FFFFD00000;
            9'h15a: data <= 64'h0000155555540000;
            9'h15b: data <= 64'h00005FFFFFF50000;
            9'h15c: data <= 64'h00007FFFFFFD0000;
            9'h15d: data <= 64'h0000555555550000;
            9'h15e: data <= 64'h0000000000000000;
            9'h15f: data <= 64'h0000000000000000;
            // CODE x11 KRÓLOWA CZARNA //////////
            9'h160: data <= 64'h0000000000000000; 
            9'h161: data <= 64'h0000000000000000;
            9'h162: data <= 64'h0000000000000000;
            9'h163: data <= 64'h0000000000000000;
            9'h164: data <= 64'h0000000000000000;
            9'h165: data <= 64'h0000000000000000;
            9'h166: data <= 64'h0000000000000000;
            9'h167: data <= 64'h0000000000000000;
            9'h168: data <= 64'h0000000000000000;
            9'h169: data <= 64'h0000000000000000;
            9'h16a: data <= 64'h0000000000000000;
            9'h16b: data <= 64'h0000000000000000;
            9'h16c: data <= 64'h0001400140014000;
            9'h16d: data <= 64'h0001D007D0074000;
            9'h16e: data <= 64'h0001F407D01F4000;
            9'h16f: data <= 64'h0001FD01407F4000;
            9'h170: data <= 64'h0001FD07D07F4000;
            9'h171: data <= 64'h0001FF5FF5FF4000;
            9'h172: data <= 64'h0001FFFFFFFF4000;
            9'h173: data <= 64'h0001FFFFFFFF4000;
            9'h174: data <= 64'h00007FFFFFFD0000;
            9'h175: data <= 64'h00001FFFFFF40000;
            9'h176: data <= 64'h0000055555500000;
            9'h177: data <= 64'h000007FFFFD00000;
            9'h178: data <= 64'h000001FFFF400000;
            9'h179: data <= 64'h0000155555540000;
            9'h17a: data <= 64'h00001FFFFFF40000;
            9'h17b: data <= 64'h0000555555550000;
            9'h17c: data <= 64'h00007FFFFFFD0000;
            9'h17d: data <= 64'h0000555555550000;
            9'h17e: data <= 64'h0000000000000000;
            9'h17f: data <= 64'h0000000000000000;
            // CODE x12 KRÓL CZARNY /////////////
            9'h180: data <= 64'h0000000000000000; 
            9'h181: data <= 64'h0000000000000000;
            9'h182: data <= 64'h0000000000000000;
            9'h183: data <= 64'h0000000000000000;
            9'h184: data <= 64'h0000000000000000;
            9'h185: data <= 64'h0000000000000000;
            9'h186: data <= 64'h0000000000000000;
            9'h187: data <= 64'h0000000140000000;
            9'h188: data <= 64'h00000007D0000000;
            9'h189: data <= 64'h00000017D4000000;
            9'h18a: data <= 64'h0000007FFD000000;
            9'h18b: data <= 64'h0000007FFD000000;
            9'h18c: data <= 64'h00000017D4000000;
            9'h18d: data <= 64'h00005507D0550000;
            9'h18e: data <= 64'h0001FF57D5FF4000;
            9'h18f: data <= 64'h0007FFF7DFFFD000;
            9'h190: data <= 64'h0007FFFD7FFFD000;
            9'h191: data <= 64'h0007FFFD7FFFD000;
            9'h192: data <= 64'h0007FFFFFFFFD000;
            9'h193: data <= 64'h0007FFFFFFFFD000;
            9'h194: data <= 64'h0007FFFFFFFFD000;
            9'h195: data <= 64'h0007FFFFFFFFD000;
            9'h196: data <= 64'h0001FFFFFFFF4000;
            9'h197: data <= 64'h0001FFFFFFFF4000;
            9'h198: data <= 64'h00007FFFFFFD0000;
            9'h199: data <= 64'h0000155555540000;
            9'h19a: data <= 64'h00001FFFFFF40000;
            9'h19b: data <= 64'h0000555555550000;
            9'h19c: data <= 64'h00007FFFFFFD0000;
            9'h19d: data <= 64'h0000555555550000;
            9'h19e: data <= 64'h0000000000000000;
            9'h19f: data <= 64'h0000000000000000;
            // CODE x13 possible move ///////////
            9'h1a0: data <= 64'h0000000000000000;   
            9'h1a1: data <= 64'h0000000000000000;
            9'h1a2: data <= 64'h0000000000000000;
            9'h1a3: data <= 64'h0000000000000000;
            9'h1a4: data <= 64'h0000000000000000;
            9'h1a5: data <= 64'h0000000000000000;
            9'h1a6: data <= 64'h0000000000000000;
            9'h1a7: data <= 64'h0000000000000000;
            9'h1a8: data <= 64'h0000000000000000;
            9'h1a9: data <= 64'h0000000000000000;
            9'h1aa: data <= 64'h0000000000000000;
            9'h1ab: data <= 64'h0000000000000000; 
            9'h1ac: data <= 64'h0000000550000000; 
            9'h1ad: data <= 64'h0000001554000000; 
            9'h1ae: data <= 64'h0000005555000000; 
            9'h1af: data <= 64'h0000005555000000;
            9'h1b0: data <= 64'h0000005555000000;
            9'h1b1: data <= 64'h0000005555000000;
            9'h1b2: data <= 64'h0000001554000000;
            9'h1b3: data <= 64'h0000000550000000;
            9'h1b4: data <= 64'h0000000000000000;
            9'h1b5: data <= 64'h0000000000000000;
            9'h1b6: data <= 64'h0000000000000000;
            9'h1b7: data <= 64'h0000000000000000;
            9'h1b8: data <= 64'h0000000000000000;
            9'h1b9: data <= 64'h0000000000000000;
            9'h1ba: data <= 64'h0000000000000000;
            9'h1bb: data <= 64'h0000000000000000;
            9'h1bc: data <= 64'h0000000000000000;
            9'h1bd: data <= 64'h0000000000000000;
            9'h1be: data <= 64'h0000000000000000;
            9'h1bf: data <= 64'h0000000000000000;
        endcase
        figure_line_pixels <= data;
    end
endmodule
